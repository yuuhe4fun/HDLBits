// module my_dff8 ( input clk, input [7:0] d, output [7:0] q );

module top_module ( 
    input clk, 
    input [7:0] d, 
    input [1:0] sel, 
    output [7:0] q 
);
    
endmodule
