// module my_dff ( input clk, input d, output q );

module top_module ( input clk, input d, output q );

    
endmodule
