module top_module (
    output out);

    assign out = 1'b0;
endmodule

// Warning (13024): Output pins are stuck at VCC or GND