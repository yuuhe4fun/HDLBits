module top_module (
    input clk,
    input d, 
    input ar,   // asynchronous reset
    output q);

endmodule
