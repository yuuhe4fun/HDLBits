module top_module (
    input clk,
    input x,
    output z
); 
    reg q1, q2, q3;
    parameter q1 = 1'b0,
              q2 = 1'b0,
              q3 = 1'b0,;
endmodule
