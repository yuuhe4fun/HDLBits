module top_module( 
    input [99:0] a, b,
    input cin,
    output [99:0] cout,
    output [99:0] sum );

    integer j;

    always @(*) begin
        for (j = 0; j <= 99; j = j + 1) begin
            
        end
    end
endmodule
